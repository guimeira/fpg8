`timescale 1ns / 1ps

module memory_controller(
	//Device clock:
	input clk,
	//Reset signal:
	input rst,
	//Signals to interface with this controller:
	//When HIGH, performs a read:
	input read,
	//When HIGH, performs a write (highest precedence over read):
	input write,
	//Address to read or write:
	input[25:0] address,
	//Data to be written:
	input[15:0] write_data,
	//Read data:
	output[15:0] read_data,
	//When high indicates that an operation is being performed:
	output busy,
	
	//Signals generated by the controller to drive the memory:
	//Memory address bus:
	output reg[25:0] mem_address,
	//Memory output enable:
	output mem_oe,
	//Memory write enable:
	output mem_we,
	//Memory clock:
	output mem_clk,
	//Memory address valid:
	output mem_adv,
	//Memory chip enable:
	output mem_mt_ce,
	//Memory upper byte:
	output mem_mt_ub,
	//Memory lower byte:
	output mem_mt_lb,
	//Memory control register enable:
	output mem_mt_cre,
	//Flash chip enable (used to disable FLASH chip):
	output flash_ce,
	//Memory data bus:
	inout[15:0] data
);
	//State machine states:
	parameter[1:0] STATE_IDLE = 2'd0, STATE_READING = 2'd1, STATE_WRITING = 2'd2;
	reg[1:0] current_state, next_state;
	
	//This ALWAYS statement controls the state transition for the state machine:
	always @(posedge clk, posedge rst) begin
		if(rst)
			current_state <= STATE_IDLE;
		else
			current_state <= next_state;
	end
	
	//This ALWAYS statement is combinational and generates the next state for the
	//state machine. The state transition is simple, when the WRITE or the READ signals
	//are HIGH, the machine goes to the appropriate state, which starts a counter.
	//When the counter reaches 6 the reading or writing cycle is over and the machine
	//returns to IDLE state. The rest of the logic in this module is derived from the current
	//state of this machine:
	always @(current_state,read,write,counter) begin
		//Set this value to avoid latches:
		next_state = current_state;
		
		case(current_state)
			STATE_IDLE: begin
				if(write) begin
					next_state = STATE_WRITING;
				end
				else if(read) begin
					next_state = STATE_READING;
				end
				else begin
					next_state = current_state;
				end
			end
			STATE_WRITING: begin
				if(counter == 3'd6) begin
					next_state = STATE_IDLE;
				end
				else begin
					next_state = STATE_WRITING;
				end
			end
			STATE_READING: begin
				if(counter == 3'd6) begin
					next_state = STATE_IDLE;
				end
				else begin
					next_state = STATE_READING;
				end
			end
		endcase
	end
	
	//This ALWAYS statement controls the address bus.
	//When we want to perform a read or write the address is copied to a register
	//so that the module that is using this controller does not need to hold the
	//address value (for whatever reason it doesnt want to).
	always @(posedge clk, posedge rst) begin
		if(rst)
			mem_address <= 26'd0;
		else begin
			if(current_state == STATE_IDLE && (read || write))
				mem_address <= address;
			else
				mem_address <= mem_address;
		end
	end
	
	//This counter is used for the timing. A reading or writing cycle is 70ns long.
	//As this module is clocked at 100MHz, each clock cycle is 10ns long, so we need
	//to count from 0 to 6 to make sure the timing requirement is fulfilled.
	reg[2:0] counter;
	always @(posedge clk, posedge rst) begin
		if(rst)
			counter <= 3'd0;
		else begin
			if(current_state != STATE_IDLE)
				counter <= counter + 3'd1;
			else
				counter <= 3'd0;
		end
	end
	
	//When writing, this register will store the data to be stored, so that the module
	//that is using this controller does not need to hold that value.
	//When reading, this register will hold the value that the memory puts on the data bus
	//after the reading cycle is finished, so that it can be accessed later.
	reg[15:0] data_reg;
	always @(posedge clk, posedge rst) begin
		if(rst)
			data_reg <= 16'd0;
		else begin
			if(current_state == STATE_IDLE && write)
				data_reg <= write_data;
			else if(current_state == STATE_READING && counter == 3'd6)
				data_reg <= data;
			else
				data_reg <= data_reg;
		end
	end
	
	//The data read from the memory:
	assign read_data = data_reg;
	
	//Tri-state on data bus:
	assign data = current_state == STATE_WRITING ? data_reg : 16'bzzzzzzzzzzzzzzzz;
	
	//Busy is high whenever we are not in STATE_IDLE:
	assign busy = current_state != STATE_IDLE;
	
	//Output enable is LOW when we are in STATE_READING:
	assign mem_oe = current_state != STATE_READING;
	
	//Write enable is LOW when we are in STATE_WRITING:
	assign mem_we = current_state != STATE_WRITING;
	
	//The memory clock is always on LOW for asynchronous mode:
	assign mem_clk = 1'b0;
	
	//The address valid signal is always on LOW for asynchronous mode:
	assign mem_adv = 1'b0;
	
	//The chip enable signal is LOW to enable the memory chip:
	assign mem_mt_ce = 1'b0;
	
	//Activate the upper byte:
	assign mem_mt_ub = 1'b0;
	
	//Activate the lower byte:
	assign mem_mt_lb = 1'b0;
	
	//The chip register is not used in asynchronous mode:
	assign mem_mt_cre = 1'b0;
	
	//Disable the FLASH chip:
	assign flash_ce = 1'b1;
endmodule
